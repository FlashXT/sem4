<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-29.5792,4.19583,74.9708,-47.8542</PageViewport>
<gate>
<ID>2</ID>
<type>AE_OR4</type>
<position>53.5,-30</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>21 </input>
<input>
<ID>IN_3</ID>22 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND3</type>
<position>38.5,-20.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>24 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND3</type>
<position>38.5,-27</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>25 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND3</type>
<position>38.5,-33.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<input>
<ID>IN_2</ID>26 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND3</type>
<position>38.5,-40</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>32 </input>
<input>
<ID>IN_2</ID>27 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>25,-22.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>25,-29</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>25,-35.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>25,-42</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>30,-7</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>33,-7</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_SMALL_INVERTER</type>
<position>31.5,-14</position>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_SMALL_INVERTER</type>
<position>34.5,-14</position>
<input>
<ID>IN_0</ID>31 </input>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>-1,-32.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>-1.5,-39</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_OR2</type>
<position>7,-35.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_SMALL_INVERTER</type>
<position>-12,-35</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>-7.5,-40</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>-7,-33.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>-12,-28.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_MUX_2x1</type>
<position>-13.5,-14.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>4 </output>
<input>
<ID>SEL_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>-18,-15.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>-18,-13.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>-13.5,-9.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>59.5,-30</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>-10,-14.5</position>
<input>
<ID>N_in0</ID>4 </input>
<input>
<ID>N_in3</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>12,-35.5</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AE_MUX_4x1</type>
<position>10,-15</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>7 </input>
<output>
<ID>OUT</ID>11 </output>
<input>
<ID>SEL_0</ID>6 </input>
<input>
<ID>SEL_1</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>3.5,-11</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>3.5,-16</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>3.5,-18.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>3.5,-13.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>10,-7</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>12,-7</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>15,-15</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>57,1</position>
<gparam>LABEL_TEXT SAMARTH KOSTA</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>-7.5,-14</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>17.5,-14.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>-20.5,-13.5</position>
<gparam>LABEL_TEXT 11</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>-20.5,-15.5</position>
<gparam>LABEL_TEXT 10</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>14.5,-35</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>-10,-39.5</position>
<gparam>LABEL_TEXT 11</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>-9.5,-33.5</position>
<gparam>LABEL_TEXT 10</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>22.5,-42</position>
<gparam>LABEL_TEXT 10</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>22.5,-35.5</position>
<gparam>LABEL_TEXT 11</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>22.5,-29</position>
<gparam>LABEL_TEXT 12</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>22.5,-22.5</position>
<gparam>LABEL_TEXT 13</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>29,-4</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>33.5,-4</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>63,-29.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>-12,-26</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>-13.5,-7</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>13,-4.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>9,-4.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-12,-13.5,-11.5</points>
<connection>
<GID>33</GID>
<name>SEL_0</name></connection>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16,-13.5,-15.5,-13.5</points>
<connection>
<GID>33</GID>
<name>IN_1</name></connection>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-16,-15.5,-15.5,-15.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-14.5,-9,-14.5</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>N_in0</name></connection>
<intersection>-9 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-9,-14.5,-9,-13.5</points>
<intersection>-14.5 1</intersection>
<intersection>-13.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-10,-13.5,-9,-13.5</points>
<connection>
<GID>40</GID>
<name>N_in3</name></connection>
<intersection>-9 3</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-10,10,-9</points>
<connection>
<GID>44</GID>
<name>SEL_1</name></connection>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-10,11,-9.5</points>
<connection>
<GID>44</GID>
<name>SEL_0</name></connection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11,-9.5,12,-9.5</points>
<intersection>11 0</intersection>
<intersection>12 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12,-9.5,12,-9</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-12,6.5,-11</points>
<intersection>-12 3</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-11,6.5,-11</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>6.5,-12,7,-12</points>
<connection>
<GID>44</GID>
<name>IN_3</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-14,7,-14</points>
<connection>
<GID>44</GID>
<name>IN_2</name></connection>
<intersection>6 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>6,-14,6,-13.5</points>
<intersection>-14 1</intersection>
<intersection>-13.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>5.5,-13.5,6,-13.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>6 3</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-16,7,-16</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>6.5,-18,7,-18</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>6.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>6.5,-18.5,6.5,-18</points>
<intersection>-18.5 5</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>5.5,-18.5,6.5,-18.5</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>6.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-15,14,-15</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<connection>
<GID>52</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-35.5,11,-35.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<connection>
<GID>42</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2,-32.5,3,-32.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>3 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>3,-34.5,3,-32.5</points>
<intersection>-34.5 6</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>3,-34.5,4,-34.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>3 4</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-39,3,-36.5</points>
<intersection>-39 2</intersection>
<intersection>-36.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>1.5,-39,3,-39</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>3,-36.5,4,-36.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-40,-4.5,-40</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5,-33.5,-4,-33.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-33,-12,-30.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>-31.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-12,-31.5,-4,-31.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-38,-12,-37</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,-38,-4.5,-38</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-27,47.5,-20.5</points>
<intersection>-27 1</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-27,50.5,-27</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-20.5,47.5,-20.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-29,46,-27</points>
<intersection>-29 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-29,50.5,-29</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-27,46,-27</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-33.5,46,-31</points>
<intersection>-33.5 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-31,50.5,-31</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-33.5,46,-33.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-40,47.5,-33</points>
<intersection>-40 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-33,50.5,-33</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-40,47.5,-40</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-30,58.5,-30</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>38</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-22.5,35.5,-22.5</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-29,35.5,-29</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-35.5,35.5,-35.5</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-42,35.5,-42</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-27,30,-9</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>-27 6</intersection>
<intersection>-20.5 9</intersection>
<intersection>-12 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>30,-27,35.5,-27</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>30,-12,31.5,-12</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>30,-20.5,35.5,-20.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-31.5,33,-9</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>-31.5 9</intersection>
<intersection>-18.5 8</intersection>
<intersection>-12 11</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>33,-18.5,35.5,-18.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>33,-31.5,35.5,-31.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>33,-12,34.5,-12</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-40,31.5,-16</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>-40 1</intersection>
<intersection>-33.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-40,35.5,-40</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-33.5,35.5,-33.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-38,34.5,-16</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-38 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-38,35.5,-38</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-25,35.5,-25</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 9></circuit>