<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0.624998,-4.525,79.0375,-43.5625</PageViewport>
<gate>
<ID>2</ID>
<type>AI_XOR2</type>
<position>12,-36</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>12,-40.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>17.5,-36</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>17.5,-40.5</position>
<input>
<ID>N_in0</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>8,-30.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>5,-30.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>22.5,-35.5</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>42,-31.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_AND2</type>
<position>42,-36</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>42,-40.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_OR3</type>
<position>50.5,-36</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>7 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>22</ID>
<type>AI_XOR2</type>
<position>50.5,-24</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AI_XOR2</type>
<position>42,-20</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>57.5,-24</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>GA_LED</type>
<position>57.5,-36</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>37.5,-14</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>35,-14</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>32.5,-14</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>66.5,-5.5</position>
<gparam>LABEL_TEXT SAMARTH KOSTA</gparam>
<gparam>TEXT_HEIGHT 1.7</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>24,-40</position>
<gparam>LABEL_TEXT CARRY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>5,-27</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>8,-27</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>12,-23.5</position>
<gparam>LABEL_TEXT HALF ADDER</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>38,-7.5</position>
<gparam>LABEL_TEXT FULL ADDER</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>32.5,-11</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>35,-11</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>37.5,-11</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>63,-23.5</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>65,-35.5</position>
<gparam>LABEL_TEXT CARRY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-40.5,16.5,-40.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-36,16.5,-36</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>6</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-41.5,5,-32.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-41.5 1</intersection>
<intersection>-37 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-41.5,9,-41.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>5,-37,9,-37</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-39.5,8,-32.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 3</intersection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-35,9,-35</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>8,-39.5,9,-39.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-24,56.5,-24</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<connection>
<GID>24</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-36,56.5,-36</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<connection>
<GID>25</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-40.5,46,-38</points>
<intersection>-40.5 2</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-38,47.5,-38</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-40.5,46,-40.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-36,47.5,-36</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-34,46,-31.5</points>
<intersection>-34 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-34,47.5,-34</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-31.5,46,-31.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-23,46,-20</points>
<intersection>-23 1</intersection>
<intersection>-20 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-23,47.5,-23</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>45,-20,46,-20</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-41.5,32.5,-16</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-41.5 1</intersection>
<intersection>-37 5</intersection>
<intersection>-25 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-41.5,39,-41.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32.5,-25,47.5,-25</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>32.5,-37,39,-37</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-39.5,37.5,-16</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 1</intersection>
<intersection>-30.5 2</intersection>
<intersection>-19 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-39.5,39,-39.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-30.5,39,-30.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>37.5,-19,39,-19</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-35,35,-16</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>-35 1</intersection>
<intersection>-32.5 3</intersection>
<intersection>-21 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-35,39,-35</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-32.5,39,-32.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>35,-21,39,-21</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 9></circuit>