<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>8.35,2.875,112.9,-49.175</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>33.5,-29</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AI_XOR2</type>
<position>33.5,-24</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_SMALL_INVERTER</type>
<position>27.5,-30</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>38.5,-24</position>
<input>
<ID>N_in0</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>38.5,-29</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>27.5,-19.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>24.5,-19.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>24.5,-16.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>27.5,-16.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>44.5,-23.5</position>
<gparam>LABEL_TEXT D = A-B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>43,-28.5</position>
<gparam>LABEL_TEXT Bout</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>64,-14</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>61,-14</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>61,-11</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>64,-11</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>67,-14</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>67,-11</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_AND2</type>
<position>76,-30.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_AND2</type>
<position>76,-35.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND2</type>
<position>76,-40.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_OR3</type>
<position>84,-35.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>89,-35.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AE_SMALL_INVERTER</type>
<position>70,-39.5</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_SMALL_INVERTER</type>
<position>70,-31.5</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AO_XNOR2</type>
<position>84,-23</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>AO_XNOR2</type>
<position>76,-20</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>89,-23</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>95,-22.5</position>
<gparam>LABEL_TEXT D = A-B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>93.5,-35</position>
<gparam>LABEL_TEXT Bout</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>29.5,-7</position>
<gparam>LABEL_TEXT HALF SUBTRACTOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>76,-7</position>
<gparam>LABEL_TEXT FULL SUBTRACTOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>98,1.5</position>
<gparam>LABEL_TEXT SAMARTH KOSTA</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>36.5,-24,37.5,-24</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>36.5,-29,37.5,-29</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>10</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-30,30.5,-30</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-28,27.5,-21.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-28 3</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-23,30.5,-23</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27.5,-28,30.5,-28</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-30,24.5,-21.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-30 1</intersection>
<intersection>-25 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-30,25.5,-30</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24.5,-25,30.5,-25</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>10</ID>
<points>79,-35.5,81,-35.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<connection>
<GID>31</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-33.5,80,-30.5</points>
<intersection>-33.5 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-33.5,81,-33.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79,-30.5,80,-30.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-40.5,80,-37.5</points>
<intersection>-40.5 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-37.5,81,-37.5</points>
<connection>
<GID>31</GID>
<name>IN_2</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79,-40.5,80,-40.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87,-35.5,88,-35.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<connection>
<GID>32</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-31.5,73,-31.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-39.5,73,-39.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-41.5,64,-16</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-41.5 1</intersection>
<intersection>-34.5 3</intersection>
<intersection>-21 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-41.5,73,-41.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,-34.5,73,-34.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>64,-21,73,-21</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-39.5,61,-16</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 1</intersection>
<intersection>-31.5 3</intersection>
<intersection>-19 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-39.5,68,-39.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>61,-31.5,68,-31.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>61,-19,73,-19</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-36.5,67,-16</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-36.5 1</intersection>
<intersection>-29.5 3</intersection>
<intersection>-24 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-36.5,73,-36.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>67,-29.5,73,-29.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>67,-24,81,-24</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79,-20,80,-20</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>80 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>80,-22,80,-20</points>
<intersection>-22 10</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>80,-22,81,-22</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>80 9</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87,-23,88,-23</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-69.4</PageViewport></page 9></circuit>